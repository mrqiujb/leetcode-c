module s9234(clock);

input wire clock;

endmodule

